// INSTRUCTION MEMORY

module imem #(parameter N=32)
			 (input logic [6:0] addr,
			  output logic [N-1:0] q);

	logic [N-1:0] ROM [0:127];
	
	initial
	begin	
ROM [0:59] ='{
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h8b030041,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h8b010062, //exc vector
32'h8b0600a4,
32'hd61f0200,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000
};


	end
	
	assign q = ROM[addr];
endmodule
